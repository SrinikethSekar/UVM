interface d_int;
  logic   clk;
  logic   rst;
  logic     d;
  logic     q;
  logic   q_b;
  
endinterface
